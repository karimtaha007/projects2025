module ALI_with_control();


endmodule

