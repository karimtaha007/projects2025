library verilog;
use verilog.vl_types.all;
entity orag_v2_vlg_vec_tst is
end orag_v2_vlg_vec_tst;
