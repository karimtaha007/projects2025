library verilog;
use verilog.vl_types.all;
entity arthimtic_circuit_vlg_vec_tst is
end arthimtic_circuit_vlg_vec_tst;
