library verilog;
use verilog.vl_types.all;
entity T_reg_vlg_vec_tst is
end T_reg_vlg_vec_tst;
