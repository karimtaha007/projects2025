library verilog;
use verilog.vl_types.all;
entity reg_8_bit_vlg_vec_tst is
end reg_8_bit_vlg_vec_tst;
