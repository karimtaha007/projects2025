library verilog;
use verilog.vl_types.all;
entity Memory16X10_vlg_vec_tst is
end Memory16X10_vlg_vec_tst;
