library verilog;
use verilog.vl_types.all;
entity state_controller_vlg_vec_tst is
end state_controller_vlg_vec_tst;
