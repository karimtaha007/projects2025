module reg_8_bit (output Q8,output [7:0] Q ,input [7:0] data ,input sign,load,clk,reset) ;


one_bit_reg r0(Q[0],data[0],load,clk,reset),
				r1(Q[1],data[1],load,clk,reset),
				r2(Q[2],data[2],load,clk,reset),
				r3(Q[3],data[3],load,clk,reset),
				r4(Q[4],data[4],load,clk,reset),
				r5(Q[5],data[5],load,clk,reset),
				r6(Q[6],data[6],load,clk,reset),
				r7(Q[7],data[7],load,clk,reset);
				assign Q8 =sign  ;

endmodule 