library verilog;
use verilog.vl_types.all;
entity one_bit_reg_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end one_bit_reg_vlg_check_tst;
