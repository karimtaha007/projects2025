library verilog;
use verilog.vl_types.all;
entity control_unit_test_vlg_vec_tst is
end control_unit_test_vlg_vec_tst;
