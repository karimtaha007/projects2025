library verilog;
use verilog.vl_types.all;
entity logic_circuit_vlg_vec_tst is
end logic_circuit_vlg_vec_tst;
