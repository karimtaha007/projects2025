library verilog;
use verilog.vl_types.all;
entity one_bit_reg_vlg_vec_tst is
end one_bit_reg_vlg_vec_tst;
