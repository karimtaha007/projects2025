library verilog;
use verilog.vl_types.all;
entity mux4x1_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux4x1_vlg_check_tst;
