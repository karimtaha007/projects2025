Smodule D_FF (output reg Q , input D,clk,reset ) ; 

always @(posedge clk )
begin
if(reset == 1) 
	Q <= 1'b0 ; 
else 
	Q <=  D ; 

end 



endmodule